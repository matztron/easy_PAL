module OR_MATRIX (
    //
);


endmodule